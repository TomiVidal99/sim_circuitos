* La idea de este script es automatizar la simulación de variación de parámetros
* Se ajustan los valores de resistencias, Capacitancias e Inductancias que se van a emplear
* Y luego en el circuito se reemplaza de la siguiente manera:
*
* Si quiero una resistencia al 10% y evaluar el peor caso cuando es más grande, es decir 1.1 veces su valor se usa:
* {R1_10_}
*
* En cambio si quiero evaluar la misma resistencia cuando es el peor caso cuando vale lo menos posible:
* {R1_10}
*
* Y así de fácil se pueden evaluar diferentes valores, en vez de estar calculándolos a mano.
*
* POR AHORA SOLO HAY AL 10%, 5% y 1%. PERO SE PUEDE EXTENDER FACILMENTE

* Resistencias
.param R1=10k
.param R2=10k
.param R3=10k
.param R4=10k
.param R5=10k
.param R6=10k
.param R7=10k
.param R8=10k
.param R9=10k
.param R10=10k
.param R11=10k
.param R12=10k
.param R13=10k
.param R14=10k
.param R15=10k
.param R16=10k
.param R17=10k
.param R18=10k
.param R19=10k
.param R20=10k

* Capacitancias
.param C1=100u
.param C2=100u
.param C3=100u
.param C4=100u
.param C5=100u
.param C6=100u
.param C7=100u
.param C8=100u
.param C9=100u
.param C10=100u
.param C11=100u
.param C12=100u
.param C13=100u
.param C14=100u
.param C15=100u
.param C16=100u
.param C17=100u
.param C18=100u
.param C19=100u
.param C20=100u

* Inductancias
.param L1=100u
.param L2=100u
.param L3=100u
.param L4=100u
.param L5=100u
.param L6=100u
.param L7=100u
.param L8=100u
.param L9=100u
.param L10=100u
.param L11=100u
.param L12=100u
.param L13=100u
.param L14=100u
.param L15=100u
.param L16=100u
.param L17=100u
.param L18=100u
.param L19=100u
.param L20=100u
* ---------------------------

* ---------------- Resistencias ----------------
.param R1_10_=R1*0.9
.param R2_10_=R2*0.9
.param R3_10_=R3*0.9
.param R4_10_=R4*0.9
.param R5_10_=R5*0.9
.param R6_10_=R6*0.9
.param R7_10_=R7*0.9
.param R8_10_=R8*0.9
.param R9_10_=R9*0.9
.param R10_10_=R10*0.9
.param R11_10_=R11*0.9
.param R12_10_=R12*0.9
.param R13_10_=R13*0.9
.param R14_10_=R14*0.9
.param R15_10_=R15*0.9
.param R16_10_=R16*0.9
.param R17_10_=R17*0.9
.param R18_10_=R18*0.9
.param R19_10_=R19*0.9
.param R20_10_=R20*0.9

.param R1_10_=R1*1.1
.param R2_10_=R2*1.1
.param R3_10_=R3*1.1
.param R4_10_=R4*1.1
.param R5_10_=R5*1.1
.param R6_10_=R6*1.1
.param R7_10_=R7*1.1
.param R8_10_=R8*1.1
.param R9_10_=R9*1.1
.param R10_10_=R10*1.1
.param R11_10_=R11*1.1
.param R12_10_=R12*1.1
.param R13_10_=R13*1.1
.param R14_10_=R14*1.1
.param R15_10_=R15*1.1
.param R16_10_=R16*1.1
.param R17_10_=R17*1.1
.param R18_10_=R18*1.1
.param R19_10_=R19*1.1
.param R20_10_=R20*1.1

.param R1_5_=R1*0.95
.param R2_5_=R2*0.95
.param R3_5_=R3*0.95
.param R4_5_=R4*0.95
.param R5_5_=R5*0.95
.param R6_5_=R6*0.95
.param R7_5_=R7*0.95
.param R8_5_=R8*0.95
.param R9_5_=R9*0.95
.param R10_5_=R10*0.95
.param R11_5_=R11*0.95
.param R12_5_=R12*0.95
.param R13_5_=R13*0.95
.param R14_5_=R14*0.95
.param R15_5_=R15*0.95
.param R16_5_=R16*0.95
.param R17_5_=R17*0.95
.param R18_5_=R18*0.95
.param R19_5_=R19*0.95
.param R20_5_=R20*0.95

.param R1_5_=R1*1.05
.param R2_5_=R2*1.05
.param R3_5_=R3*1.05
.param R4_5_=R4*1.05
.param R5_5_=R5*1.05
.param R6_5_=R6*1.05
.param R7_5_=R7*1.05
.param R8_5_=R8*1.05
.param R9_5_=R9*1.05
.param R10_5_=R10*1.05
.param R11_5_=R11*1.05
.param R12_5_=R12*1.05
.param R13_5_=R13*1.05
.param R14_5_=R14*1.05
.param R15_5_=R15*1.05
.param R16_5_=R16*1.05
.param R17_5_=R17*1.05
.param R18_5_=R18*1.05
.param R19_5_=R19*1.05
.param R20_5_=R20*1.05

.param R1_1_=R1*0.99
.param R2_1_=R2*0.99
.param R3_1_=R3*0.99
.param R4_1_=R4*0.99
.param R5_1_=R5*0.99
.param R6_1_=R6*0.99
.param R7_1_=R7*0.99
.param R8_1_=R8*0.99
.param R9_1_=R9*0.99
.param R10_1_=R10*0.99
.param R11_1_=R11*0.99
.param R12_1_=R12*0.99
.param R13_1_=R13*0.99
.param R14_1_=R14*0.99
.param R15_1_=R15*0.99
.param R16_1_=R16*0.99
.param R17_1_=R17*0.99
.param R18_1_=R18*0.99
.param R19_1_=R19*0.99
.param R20_1_=R20*0.99

.param R1_1_=R1*1.01
.param R2_1_=R2*1.01
.param R3_1_=R3*1.01
.param R4_1_=R4*1.01
.param R5_1_=R5*1.01
.param R6_1_=R6*1.01
.param R7_1_=R7*1.01
.param R8_1_=R8*1.01
.param R9_1_=R9*1.01
.param R10_1_=R10*1.01
.param R11_1_=R11*1.01
.param R12_1_=R12*1.01
.param R13_1_=R13*1.01
.param R14_1_=R14*1.01
.param R15_1_=R15*1.01
.param R16_1_=R16*1.01
.param R17_1_=R17*1.01
.param R18_1_=R18*1.01
.param R19_1_=R19*1.01
.param R20_1_=R20*1.01

* ---------------- Capacitancias ----------------
.param C1_10_=C1*0.9
.param C2_10_=C2*0.9
.param C3_10_=C3*0.9
.param C4_10_=C4*0.9
.param C5_10_=C5*0.9
.param C6_10_=C6*0.9
.param C7_10_=C7*0.9
.param C8_10_=C8*0.9
.param C9_10_=C9*0.9
.param C10_10_=C10*0.9
.param C11_10_=C11*0.9
.param C12_10_=C12*0.9
.param C13_10_=C13*0.9
.param C14_10_=C14*0.9
.param C15_10_=C15*0.9
.param C16_10_=C16*0.9
.param C17_10_=C17*0.9
.param C18_10_=C18*0.9
.param C19_10_=C19*0.9
.param C20_10_=C20*0.9

.param C1_10_=C1*1.1
.param C2_10_=C2*1.1
.param C3_10_=C3*1.1
.param C4_10_=C4*1.1
.param C5_10_=C5*1.1
.param C6_10_=C6*1.1
.param C7_10_=C7*1.1
.param C8_10_=C8*1.1
.param C9_10_=C9*1.1
.param C10_10_=C10*1.1
.param C11_10_=C11*1.1
.param C12_10_=C12*1.1
.param C13_10_=C13*1.1
.param C14_10_=C14*1.1
.param C15_10_=C15*1.1
.param C16_10_=C16*1.1
.param C17_10_=C17*1.1
.param C18_10_=C18*1.1
.param C19_10_=C19*1.1
.param C20_10_=C20*1.1

.param C1_5_=C1*0.95
.param C2_5_=C2*0.95
.param C3_5_=C3*0.95
.param C4_5_=C4*0.95
.param C5_5_=C5*0.95
.param C6_5_=C6*0.95
.param C7_5_=C7*0.95
.param C8_5_=C8*0.95
.param C9_5_=C9*0.95
.param C10_5_=C10*0.95
.param C11_5_=C11*0.95
.param C12_5_=C12*0.95
.param C13_5_=C13*0.95
.param C14_5_=C14*0.95
.param C15_5_=C15*0.95
.param C16_5_=C16*0.95
.param C17_5_=C17*0.95
.param C18_5_=C18*0.95
.param C19_5_=C19*0.95
.param C20_5_=C20*0.95

.param C1_5_=C1*1.05
.param C2_5_=C2*1.05
.param C3_5_=C3*1.05
.param C4_5_=C4*1.05
.param C5_5_=C5*1.05
.param C6_5_=C6*1.05
.param C7_5_=C7*1.05
.param C8_5_=C8*1.05
.param C9_5_=C9*1.05
.param C10_5_=C10*1.05
.param C11_5_=C11*1.05
.param C12_5_=C12*1.05
.param C13_5_=C13*1.05
.param C14_5_=C14*1.05
.param C15_5_=C15*1.05
.param C16_5_=C16*1.05
.param C17_5_=C17*1.05
.param C18_5_=C18*1.05
.param C19_5_=C19*1.05
.param C20_5_=C20*1.05

.param C1_1_=C1*0.99
.param C2_1_=C2*0.99
.param C3_1_=C3*0.99
.param C4_1_=C4*0.99
.param C5_1_=C5*0.99
.param C6_1_=C6*0.99
.param C7_1_=C7*0.99
.param C8_1_=C8*0.99
.param C9_1_=C9*0.99
.param C10_1_=C10*0.99
.param C11_1_=C11*0.99
.param C12_1_=C12*0.99
.param C13_1_=C13*0.99
.param C14_1_=C14*0.99
.param C15_1_=C15*0.99
.param C16_1_=C16*0.99
.param C17_1_=C17*0.99
.param C18_1_=C18*0.99
.param C19_1_=C19*0.99
.param C20_1_=C20*0.99

.param C1_1_=C1*1.01
.param C2_1_=C2*1.01
.param C3_1_=C3*1.01
.param C4_1_=C4*1.01
.param C5_1_=C5*1.01
.param C6_1_=C6*1.01
.param C7_1_=C7*1.01
.param C8_1_=C8*1.01
.param C9_1_=C9*1.01
.param C10_1_=C10*1.01
.param C11_1_=C11*1.01
.param C12_1_=C12*1.01
.param C13_1_=C13*1.01
.param C14_1_=C14*1.01
.param C15_1_=C15*1.01
.param C16_1_=C16*1.01
.param C17_1_=C17*1.01
.param C18_1_=C18*1.01
.param C19_1_=C19*1.01
.param C20_1_=C20*1.01

* ---------------- Inductancias ----------------
.param L1_10_=L1*0.9
.param L2_10_=L2*0.9
.param L3_10_=L3*0.9
.param L4_10_=L4*0.9
.param L5_10_=L5*0.9
.param L6_10_=L6*0.9
.param L7_10_=L7*0.9
.param L8_10_=L8*0.9
.param L9_10_=L9*0.9
.param L10_10_=L10*0.9
.param L11_10_=L11*0.9
.param L12_10_=L12*0.9
.param L13_10_=L13*0.9
.param L14_10_=L14*0.9
.param L15_10_=L15*0.9
.param L16_10_=L16*0.9
.param L17_10_=L17*0.9
.param L18_10_=L18*0.9
.param L19_10_=L19*0.9
.param L20_10_=L20*0.9

.param L1_10_=L1*1.1
.param L2_10_=L2*1.1
.param L3_10_=L3*1.1
.param L4_10_=L4*1.1
.param L5_10_=L5*1.1
.param L6_10_=L6*1.1
.param L7_10_=L7*1.1
.param L8_10_=L8*1.1
.param L9_10_=L9*1.1
.param L10_10_=L10*1.1
.param L11_10_=L11*1.1
.param L12_10_=L12*1.1
.param L13_10_=L13*1.1
.param L14_10_=L14*1.1
.param L15_10_=L15*1.1
.param L16_10_=L16*1.1
.param L17_10_=L17*1.1
.param L18_10_=L18*1.1
.param L19_10_=L19*1.1
.param L20_10_=L20*1.1

.param L1_5_=L1*0.95
.param L2_5_=L2*0.95
.param L3_5_=L3*0.95
.param L4_5_=L4*0.95
.param L5_5_=L5*0.95
.param L6_5_=L6*0.95
.param L7_5_=L7*0.95
.param L8_5_=L8*0.95
.param L9_5_=L9*0.95
.param L10_5_=L10*0.95
.param L11_5_=L11*0.95
.param L12_5_=L12*0.95
.param L13_5_=L13*0.95
.param L14_5_=L14*0.95
.param L15_5_=L15*0.95
.param L16_5_=L16*0.95
.param L17_5_=L17*0.95
.param L18_5_=L18*0.95
.param L19_5_=L19*0.95
.param L20_5_=L20*0.95

.param L1_5_=L1*1.05
.param L2_5_=L2*1.05
.param L3_5_=L3*1.05
.param L4_5_=L4*1.05
.param L5_5_=L5*1.05
.param L6_5_=L6*1.05
.param L7_5_=L7*1.05
.param L8_5_=L8*1.05
.param L9_5_=L9*1.05
.param L10_5_=L10*1.05
.param L11_5_=L11*1.05
.param L12_5_=L12*1.05
.param L13_5_=L13*1.05
.param L14_5_=L14*1.05
.param L15_5_=L15*1.05
.param L16_5_=L16*1.05
.param L17_5_=L17*1.05
.param L18_5_=L18*1.05
.param L19_5_=L19*1.05
.param L20_5_=L20*1.05

.param L1_1_=L1*0.99
.param L2_1_=L2*0.99
.param L3_1_=L3*0.99
.param L4_1_=L4*0.99
.param L5_1_=L5*0.99
.param L6_1_=L6*0.99
.param L7_1_=L7*0.99
.param L8_1_=L8*0.99
.param L9_1_=L9*0.99
.param L10_1_=L10*0.99
.param L11_1_=L11*0.99
.param L12_1_=L12*0.99
.param L13_1_=L13*0.99
.param L14_1_=L14*0.99
.param L15_1_=L15*0.99
.param L16_1_=L16*0.99
.param L17_1_=L17*0.99
.param L18_1_=L18*0.99
.param L19_1_=L19*0.99
.param L20_1_=L20*0.99

.param L1_1_=L1*1.01
.param L2_1_=L2*1.01
.param L3_1_=L3*1.01
.param L4_1_=L4*1.01
.param L5_1_=L5*1.01
.param L6_1_=L6*1.01
.param L7_1_=L7*1.01
.param L8_1_=L8*1.01
.param L9_1_=L9*1.01
.param L10_1_=L10*1.01
.param L11_1_=L11*1.01
.param L12_1_=L12*1.01
.param L13_1_=L13*1.01
.param L14_1_=L14*1.01
.param L15_1_=L15*1.01
.param L16_1_=L16*1.01
.param L17_1_=L17*1.01
.param L18_1_=L18*1.01
.param L19_1_=L19*1.01
.param L20_1_=L20*1.01